LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

PACKAGE cpu_defs_pack IS
  constant data_width       :positive :=12;   --1.1.1
  constant address_width    :positive :=12;   --1.1.2
END cpu_defs_pack;
