use subtype_package_all.all;
