package subtype_package_all is
     
       subtype mem_data in integer range 4095 downto 0;  //subtype für Spericher
       
end subtype_package_all;
