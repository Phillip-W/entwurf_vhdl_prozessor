LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE work.def_package_all.all;
ENTITY CPU IS                               -- die CPU braucht keinerlei Ports, da alles in sie integriert wird.
  
END CPU;
