LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

PACKAGE mem_defs_pack IS
  
  --Hier alle Konstanten definieren - falls nötig
  
  --Hier alle Datentypen, Subtyps definieren - falls nötig
  
  --Hier alle nötigen Funktionen angeben
  
END mem_defs_pack;
