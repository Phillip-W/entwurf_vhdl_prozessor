LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
Use work.def_package_all.all;

package mem_package_all is
  function init_memory return mem_type;      
end mem_package_all;
