-- Hier alle Subtypes als Package reinschreiben

