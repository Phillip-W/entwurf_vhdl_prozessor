PACKAGE BODY mem_defs_pack IS

  --Hier alle Funktionen definieren
  function test return opcode_type is
    begin
      return (
        0
        );
  end test;
